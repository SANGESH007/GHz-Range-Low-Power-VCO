** sch_path: /home/sangesh007/Desktop/inverter_vco.sch
**.subckt inverter_vco
vdd vdd GND 1.8
vin vin GND 1.8
XM3 vout vin GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 vout vin vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=2.745 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt



.control
	run
	set color0=white
	dc vin 0 1.8 1m
	setplot dc
	plot vout vin
	meas dc vth when vin=vout
	print vth
.endc
.save all
.end

**** end user architecture code
**.ends
.GLOBAL GND
.end
